constant ROMDATA : blocoMemoria := (
  0  => x"800012B7",
  1  => x"80028293",
  2  => x"03900313",
  3  => x"0062A023",
  4  => x"FF9FF06F",
  5  => x"00000000",
  6  => x"00000000",
  7  => x"00000000",
  8  => x"00000000",
  9  => x"00000000",
  10  => x"00000000",
  11  => x"00000000",
  12  => x"00000000",
  13  => x"00000000",
  14  => x"00000000",
  15  => x"00000000",
  16  => x"00000000",
  17  => x"00000000",
  18  => x"00000000",
  19  => x"00000000",
  20  => x"00000000",
  21  => x"00000000",
  22  => x"00000000",
  23  => x"00000000",
  24  => x"00000000",
  25  => x"00000000",
  26  => x"00000000",
  27  => x"00000000",
  28  => x"00000000",
  29  => x"00000000",
  30  => x"00000000",
  31  => x"00000000",
  32  => x"00000000",
  33  => x"00000000",
  34  => x"00000000",
  35  => x"00000000",
  36  => x"00000000",
  37  => x"00000000",
  38  => x"00000000",
  39  => x"00000000",
  40  => x"00000000",
  41  => x"00000000",
  42  => x"00000000",
  43  => x"00000000",
  44  => x"00000000",
  45  => x"00000000",
  46  => x"00000000",
  47  => x"00000000",
  48  => x"00000000",
  49  => x"00000000",
  50  => x"00000000",
  51  => x"00000000",
  52  => x"00000000",
  53  => x"00000000",
  54  => x"00000000",
  55  => x"00000000",
  56  => x"00000000",
  57  => x"00000000",
  58  => x"00000000",
  59  => x"00000000",
  60  => x"00000000",
  61  => x"00000000",
  62  => x"00000000",
  63  => x"00000000",
  64  => x"00000000",
  65  => x"00000000",
  66  => x"00000000",
  67  => x"00000000",
  68  => x"00000000",
  69  => x"00000000",
  70  => x"00000000",
  71  => x"00000000",
  72  => x"00000000",
  73  => x"00000000",
  74  => x"00000000",
  75  => x"00000000",
  76  => x"00000000",
  77  => x"00000000",
  78  => x"00000000",
  79  => x"00000000",
  80  => x"00000000",
  81  => x"00000000",
  82  => x"00000000",
  83  => x"00000000",
  84  => x"00000000",
  85  => x"00000000",
  86  => x"00000000",
  87  => x"00000000",
  88  => x"00000000",
  89  => x"00000000",
  90  => x"00000000",
  91  => x"00000000",
  92  => x"00000000",
  93  => x"00000000",
  94  => x"00000000",
  95  => x"00000000",
  96  => x"00000000",
  97  => x"00000000",
  98  => x"00000000",
  99  => x"00000000",
  100  => x"00000000",
  101  => x"00000000",
  102  => x"00000000",
  103  => x"00000000",
  104  => x"00000000",
  105  => x"00000000",
  106  => x"00000000",
  107  => x"00000000",
  108  => x"00000000",
  109  => x"00000000",
  110  => x"00000000",
  111  => x"00000000",
  112  => x"00000000",
  113  => x"00000000",
  114  => x"00000000",
  115  => x"00000000",
  116  => x"00000000",
  117  => x"00000000",
  118  => x"00000000",
  119  => x"00000000",
  120  => x"00000000",
  121  => x"00000000",
  122  => x"00000000",
  123  => x"00000000",
  124  => x"00000000",
  125  => x"00000000",
  126  => x"00000000",
  127  => x"00000000",
  128  => x"00000000",
  129  => x"00000000",
  130  => x"00000000",
  131  => x"00000000",
  132  => x"00000000",
  133  => x"00000000",
  134  => x"00000000",
  135  => x"00000000",
  136  => x"00000000",
  137  => x"00000000",
  138  => x"00000000",
  139  => x"00000000",
  140  => x"00000000",
  141  => x"00000000",
  142  => x"00000000",
  143  => x"00000000",
  144  => x"00000000",
  145  => x"00000000",
  146  => x"00000000",
  147  => x"00000000",
  148  => x"00000000",
  149  => x"00000000",
  150  => x"00000000",
  151  => x"00000000",
  152  => x"00000000",
  153  => x"00000000",
  154  => x"00000000",
  155  => x"00000000",
  156  => x"00000000",
  157  => x"00000000",
  158  => x"00000000",
  159  => x"00000000",
  160  => x"00000000",
  161  => x"00000000",
  162  => x"00000000",
  163  => x"00000000",
  164  => x"00000000",
  165  => x"00000000",
  166  => x"00000000",
  167  => x"00000000",
  168  => x"00000000",
  169  => x"00000000",
  170  => x"00000000",
  171  => x"00000000",
  172  => x"00000000",
  173  => x"00000000",
  174  => x"00000000",
  175  => x"00000000",
  176  => x"00000000",
  177  => x"00000000",
  178  => x"00000000",
  179  => x"00000000",
  180  => x"00000000",
  181  => x"00000000",
  182  => x"00000000",
  183  => x"00000000",
  184  => x"00000000",
  185  => x"00000000",
  186  => x"00000000",
  187  => x"00000000",
  188  => x"00000000",
  189  => x"00000000",
  190  => x"00000000",
  191  => x"00000000",
  192  => x"00000000",
  193  => x"00000000",
  194  => x"00000000",
  195  => x"00000000",
  196  => x"00000000",
  197  => x"00000000",
  198  => x"00000000",
  199  => x"00000000",
  200  => x"00000000",
  201  => x"00000000",
  202  => x"00000000",
  203  => x"00000000",
  204  => x"00000000",
  205  => x"00000000",
  206  => x"00000000",
  207  => x"00000000",
  208  => x"00000000",
  209  => x"00000000",
  210  => x"00000000",
  211  => x"00000000",
  212  => x"00000000",
  213  => x"00000000",
  214  => x"00000000",
  215  => x"00000000",
  216  => x"00000000",
  217  => x"00000000",
  218  => x"00000000",
  219  => x"00000000",
  220  => x"00000000",
  221  => x"00000000",
  222  => x"00000000",
  223  => x"00000000",
  224  => x"00000000",
  225  => x"00000000",
  226  => x"00000000",
  227  => x"00000000",
  228  => x"00000000",
  229  => x"00000000",
  230  => x"00000000",
  231  => x"00000000",
  232  => x"00000000",
  233  => x"00000000",
  234  => x"00000000",
  235  => x"00000000",
  236  => x"00000000",
  237  => x"00000000",
  238  => x"00000000",
  239  => x"00000000",
  240  => x"00000000",
  241  => x"00000000",
  242  => x"00000000",
  243  => x"00000000",
  244  => x"00000000",
  245  => x"00000000",
  246  => x"00000000",
  247  => x"00000000",
  248  => x"00000000",
  249  => x"00000000",
  250  => x"00000000",
  251  => x"00000000",
  252  => x"00000000",
  253  => x"00000000",
  254  => x"00000000",
  255  => x"00000000",

  -- restante zerado até 255 (se necessário ajuste memoryAddrWidth)
);

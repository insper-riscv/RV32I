constant ROMDATA : blocoMemoria := (
  0   => x"20000293",
  1   => x"00028E33",
  2   => x"00900313",
  3   => x"00030E33",
  4   => x"0062A023",
  5   => x"FF5FF06F",
  6 to 255 => x"00000000"  -- restante zerado
);
